// Module: top_hdl.sv
// Author: Rehan Iqbal
// Date: January 15th, 2018
// Organization: Portland State University
//
// Description:
//
// This module provides the top-level HDL code for Lab 1. It instantiates
// a copy of the sequence_gen module and sequence_gen_test module and
// wires them together. It also creates a 10ns clock signal to send
// to both. All control signals are generated by sequence_gen_test;
// this top-level does no simulation or hardwork work.
//
// The top-level module assumes the testbench is in a seperate directory;
// adjust the `include directive below as needed.
//
////////////////////////////////////////////////////////////////////////////////

`include "definitions.sv"
`include "../tb/sequence_gen_test_lab2.v"

module top_hdl();

	timeunit 10ns / 1ns;

	/************************************************************************/
	/* Local parameters and variables										*/
	/************************************************************************/

	ulogic1		clk	= 1'b0;

	ulogic1		reset_n;
	ulogic1		fibonacci;
	ulogic1		triangle;
	ulogic1		load;
	ulogic1		clear;
	ulogic16	order;
	ulogic64	data_in;

	ulogic1		done;
	ulogic64	data_out;
	ulogic1		overflow;
	ulogic1		error;

	/************************************************************************/
	/* Module instantiations												*/
	/************************************************************************/

	//////////////////
	// sequence_gen //
	//////////////////

	sequence_gen i_sequence_gen (

		.clk      		(clk),			// I [0] clock signal
		.reset_n  		(reset_n),		// I [0] active-low reset
		.fibonacci		(fibonacci),	// I [0] mode: perform fibonacci calculation
		.triangle 		(triangle),		// I [0] mode: perform triangle calculation
		.load     		(load),			// I [0] active (2 cycles) --> load data into FSM
		.clear    		(clear),		// I [0] clear results off 'data_out' bus
		.order    		(order),		// I [15:0] calculate the Nth value of the sequence
		.data_in  		(data_in),		// I [63:0] initial value of the sequence

		.done     		(done),			// O [0] active (1 cycle) --> data is ready
		.data_out 		(data_out),		// O [63:0] calculated value of the sequence
		.overflow 		(overflow),		// O [0] calculation exceeds bus max
		.error    		(error)			// O [0] indicates bad control input or bad data

	);

	///////////////////////
	// sequence_gen_test //
	///////////////////////

	sequence_gen_test i_sequence_gen_test (

		.clk      		(clk),			// I [0] clock signal
		.done     		(done),			// I [0] active (1 cycle) --> data is ready
		.error    		(error),		// I [0] indicates bad control input or bad data
		.overflow 		(overflow),		// I [0] calculation exceeds bus max
		.data_out 		(data_out),		// I [63:0] calculed value of the sequence

		.reset_n  		(reset_n),		// O [0] active-low reset
		.load     		(load),			// O [0] active (2 cycles) load data into FSM
		.fibonacci		(fibonacci),	// O [O] mode: perform fibonacci calculation
		.triangle 		(triangle),		// O [0] mode: perform triangle calculation
		.clear    		(clear),		// O [0] clear results off 'data_out' bus
		.order    		(order),		// O [15:0] calculate the Nth value of the sequence
		.data_in  		(data_in)		// O [63:0] initial value of the sequence

	);

	//////////////////
	// seq_gen_chkr //
	//////////////////

	seq_gen_chkr #(

		.CHKR_RULE_1	(1'b0),		// reset_n asserts -> all outputs are 0 within 1 cycle
		.CHKR_RULE_2	(1'b0),		// load asserts -> valid 'data_in' and 'order' bits
		.CHKR_RULE_3	(1'b0),		// load asserts -> either 'fibonacci' or 'triangle' active on same cycle
		.CHKR_RULE_4	(1'b0),		// done asserts -> 'data_out' correct on same cycle
		.CHKR_RULE_5	(1'b0),		// overflow asserts -> 'data_out' all 1's on same cycle
		.CHKR_RULE_6	(1'b0),		// error asserts -> 'data_out' all X's on same cycle
		.CHKR_RULE_7	(1'b0)) 	// load asserts -> 'done' and 'data_out' within <order+2> cycles

	i_seq_gen_chkr (

		.clk      		(clk),			// I [0] clock signal
		.reset_n  		(reset_n),		// I [0] active-low reset
		.fibonacci		(fibonacci),	// I [0] mode: perform fibonacci calculation
		.triangle 		(triangle),		// I [0] mode: perform triangle calculation
		.load     		(load),			// I [0] active (2 cycles) --> load data into FSM
		.clear    		(clear),		// I [0] clear results off 'data_out' bus
		.order    		(order),		// I [15:0] calculate the Nth value of the sequence
		.data_in  		(data_in),		// I [63:0] initial value of the sequence

		.done     		(done),			// I [0] active (1 cycle) --> data is ready
		.data_out 		(data_out),		// I [63:0] calculated value of the sequence
		.overflow 		(overflow),		// I [0] calculation exceeds bus max
		.error    		(error)			// I [0] indicates bad control input or bad data

	);

	/************************************************************************/
	/* initial block : clk													*/
	/************************************************************************/

	initial begin
		forever #0.5 clk = !clk;
	end

endmodule // top_hdl